module constants

pub const day_expiration_refresh_token = 2
