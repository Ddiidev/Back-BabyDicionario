module interfaces

pub interface IStorageBabydi {
	create_user(uuid string) !
}
