module models

pub enum Sexo as int {
	masculino = 0
	feminino = 1
}