module models

pub struct FamilyProfiles {
pub mut:
	father Profile
	mother Profile
	babys []Profile
}