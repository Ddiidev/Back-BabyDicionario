module constants

pub const msg_err_json_contract = 'O JSON fornecido não está de acordo com o contrato esperado.'

pub const msg_err_token_invalid = 'Token inválido'

pub const msg_err_user_not_found = 'Usuário não encontrado'

pub const msg_user_found = 'Usuário encontrado'

pub const msg_err_send_email = 'Falha ao enviar o email de confirmação'

pub const msg_err_generate_token = 'Falha ao gerar token de acesso'

pub const msg_send_email = 'Email enviado com sucesso'

pub const msg_err_not_found_email = 'Email não encontrado'

pub const msg_err_recovery_contain_recovery_password = 'Já existe uma solicitação de recuperação solicitada a pouco tempo, favor tentar novamente após 15min.'

pub const msg_err_user_fail_unblocked = 'Falha ao desbloquear a conta de usuário, por favor entre em contato com suporte via email'

pub const msg_err_email_in_use = 'Este email já foi registrado no Dicionário do bebê.\n\nPrefira fazer o login ao invés de nova conta (E pode preencher o formulário de senha esquecida caso necessário).'
