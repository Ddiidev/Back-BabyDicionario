module types

pub enum Sex {
	masculino = 0
	feminino  = 1
}
