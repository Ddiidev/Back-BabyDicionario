module contract_shared

pub enum Sex {
	masculino = 0
	feminino  = 1
}
