module constants

pub const uuid_empty = '00000000-0000-0000-0000-000000000000'
