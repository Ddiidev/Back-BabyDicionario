module entities

import contracts.profile as cprofile
import contracts.contract_shared { Sexo }
import time
import constants

@[table: 'profiles']
pub struct Profile {
pub:
	id               int        @[primary; sql: serial]
	uuid             string
	short_uuid       string
	name_shared_link string
	family_id        int
	apelido          string
	primeiro_nome    string
	segundo_nome     string
	data_nascimento  ?time.Time @[default: 'null']
	idade            f64        @[sql_type: 'NUMERIC']
	peso             f64        @[sql_type: 'NUMERIC']
	sexo             Sexo
	altura           f64        @[sql_type: 'NUMERIC']
	cor              string
	pai_id           ?int
	mae_id           ?int
	created_at       time.Time = time.utc()
	updated_at       time.Time = time.utc()
}

pub fn (p Profile) adapter() cprofile.ProfileAlias {
	return cprofile.ProfileAlias(cprofile.Profile{
		uuid: p.uuid
		apelido: p.apelido
		primeiro_nome: p.primeiro_nome
		segundo_nome: p.segundo_nome
		idade: p.idade
		peso: p.peso
		cor: p.cor
		sexo: p.sexo
		altura: p.altura
		data_nascimento: p.data_nascimento or { constants.time_empty }
	})
}

pub fn (p Profile) validated() Profile {
	return Profile{
		...p
		primeiro_nome: p.primeiro_nome.trim_space()
		segundo_nome: p.segundo_nome.trim_space()
		apelido: p.apelido.trim_space()
		cor: p.cor.trim_space()
		short_uuid: p.uuid.all_after_last('-')
		name_shared_link: p.primeiro_nome
	}
}
