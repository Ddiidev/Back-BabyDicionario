module token

pub struct TokenJwtContract {
pub:
	email string
}