module contract_shared

pub enum Sexo {
	masculino = 0
	feminino  = 1
}
