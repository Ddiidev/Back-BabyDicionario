module token

pub struct TokenContractRecoverResponse {
pub:
	access_token  string
}
