module contracts

pub type UserUUID = string