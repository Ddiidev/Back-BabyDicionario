module contract_shared

pub enum Responsible as i8 {
	pai = 0
	mae = 1
}
