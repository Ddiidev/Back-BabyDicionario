module services

import domain.profile.models

pub struct FamilyService {}

pub fn (f FamilyService) create(family models.Family) ! {
	
}