module models

pub struct TokenPayload {
pub:
	email string
}