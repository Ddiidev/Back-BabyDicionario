module interfaces

pub interface IConfig {
	get_api_storage_babydi() !string
}
