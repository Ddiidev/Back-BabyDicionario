module words

pub struct WordContract {
pub:
	profile_uuid string
	palavra      string
	traducao     string
	pronuncia    string
	audio        string
}
