module confirmation

pub struct ConfirmationEmail {
pub:
	email string
	code string
}
