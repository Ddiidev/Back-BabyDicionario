module interfaces

pub interface ITokenJwtContract {
	email string
}
