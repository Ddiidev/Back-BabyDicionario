module services

