module constants

import time

pub const time_empty = time.date_from_days_after_unix_epoch(0)
