module errors

pub struct TokenNoExist {Error}

pub struct TokenExist {Error}

pub struct RefreshTokenExpired {Error}