module constants

pub const msg_err_email_or_pass = 'Email ou senha estão incorretos.'

pub const msg_err_json_contract = 'O JSON fornecido não está de acordo com o contrato esperado.'

pub const msg_err_token_invalid = 'Token inválido'

pub const msg_err_user_not_found = 'Usuário não encontrado'

pub const msg_err_user_found = 'Usuário encontrado'