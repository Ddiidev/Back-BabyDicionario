module ws_context

import veb

pub struct Context {
	veb.Context
}
