module errors

pub struct TokenNoExist {
	Error
}

pub struct TokenAlreadyExist {
	Error
}

pub struct RefreshTokenExpired {
	Error
}
