module words

pub struct WordContract {
pub:
	profile_uuid string
}
