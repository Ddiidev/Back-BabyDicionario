module ws_context

import x.vweb

pub struct Context {
	vweb.Context
}
