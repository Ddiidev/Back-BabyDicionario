module interfaces

pub interface IToken {
	payload IPayload
	str() string
}