module interfaces

pub interface IEmailService {
	congratulations(to string, user_name string) !
}
