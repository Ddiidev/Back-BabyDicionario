module token

pub struct TokenContract {
pub:
	access_token string
	refresh_token string
}