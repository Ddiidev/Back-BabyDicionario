module confirmation

pub struct ConfirmationEmailByCode {
pub:
	email string
	code  string
}
