module tests

import net.http

fn test_contract_invalid() {
}
