module contract_shared

pub enum Responsavel as i8 {
	pai = 0
	mae = 1
}
