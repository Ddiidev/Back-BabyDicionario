module implementations

pub struct JwtRepository {}