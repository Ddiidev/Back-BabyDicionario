module types

pub type AccessToken = string