module contract_shared

pub enum Responsible as int {
	pai = 0
	mae = 1
}
