module token

// TODO: Logo se tornará obsoleto para algo que faça mais sentido
pub struct TokenJwtContract {
pub:
	email string
}
